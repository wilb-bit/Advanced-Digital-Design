module out (

);


endmodule
