module shiftReg(reset_n, loadData, dataBus, shiftClk, shiftComplete, shiftLSB);
	
	parameter bitLength = 16; // Default width
	input reset_n; // Active low reset.
	input loadData; // Active high data load.
	input [bitLength - 1:0] dataBus; // Input data bus,
	input shiftClk; // Input clock.
	
	output reg shiftComplete; // Shift complete flag
	output shiftLSB; // LSB output
	
	reg [bitLength - 1:0] shiftValue;
	reg shiftEnabled;
	integer shiftCounter;
	
	
	// Set the LSB to be output.
	assign shiftLSB = shiftValue[0];
	
	
	// Set an always block to utilise the main system clock.
	always @(posedge(shiftClk))
	begin
		// Create the reset logic
		if(reset_n == 1'b0)
			begin
				shiftValue <= 8'b00000000;
				shiftEnabled <= 1'b0;
				shiftCounter <= 0;
				shiftComplete <= 1'b0;
			end
		else if(loadData == 1'b1)
			begin
				shiftValue <= dataBus;
				shiftEnabled <= 1'b1;
				shiftCounter <= (bitLength - 1'b1);
				shiftComplete <= 1'b0;
			end
		else if ((shiftEnabled == 1'b1) && (shiftComplete == 1'b0))
			begin
				shiftValue <= shiftValue >> 1'b1;
				shiftCounter <= shiftCounter - 1'b1;
				// Check to see whether the count is complete
				if(shiftCounter == 1'b0)
				shiftComplete <= 1'b1;
			end
		else
			begin
				// Latched condition
				shiftValue <= shiftValue;
				// Check to see whether the count is complete
				if(shiftCounter == 1'b0)
				shiftComplete <= 1'b1;
			end
	end
endmodule
